���      }�(�
components�]�(}�(�element��circuit_elements��CircuitElement���)��}�(�name��I4��value�G@      �element_type��current_source��nodes�]�(K Keub�	comp_type�h�center�G@m@     G@e�     ���rotation�M�shape_points�]��	terminals�]�(J����K ��KK ��e�current_arrows�]�(MAMBe�voltage_arrows�]��current�G@      u}�(hh)��}�(h
�V10�hG@B      h�voltage_source�h]�(KK eubhh$hG@s     G@k�     ��hK h]�h]�(K J������K K��eh]�(MCMDeh]�h�numpy._core.multiarray��scalar����numpy��dtype����f8�����R�(K�<�NNNJ����J����K t�bC233333󿔆�R�u}�(hh)��}�(h
�R15�hG@(      h�resistor�h]�(KKeubhh?hG@s�     G@`@     ��hKZh]�(J����K ��J����J������K K
��K
J������KK ��eh]�(hheh]�(MEMFeh]�hh/h5C333333󿔆�R�u}�(hh)��}�(h
�R16�hG@      h�resistor�h]�(KKeubhhRhG@}@     G@W      ��hK h]�(hChDhEhFhGeh]�(hheh]�(MGMHeh]�hh/h5C������@���R�u}�(hh)��}�(h
�R17�hG@      h�resistor�h]�(KK eubhh`hG@z      G@e�     ��hKZh]�(hChDhEhFhGeh]�(hheh]�(MIMJeh]�hh/h5C������@���R�u}�(hh)��}�(h
�R18�hG@      h�resistor�h]�(KK eubhhnhG@��     G@d�     ��hKZh]�(hChDhEhFhGeh]�(hheh]�(MKMLeh]�hh/h5C������@���R�u}�(hNh�ground�hG@l�     G@t�     ��hK h]�h]�(J����K ��K
K ��e�	is_ground��h]�h]�ue�wires�]�(}�(h
�Wire1��comp1_index�K �	term1_idx�K�comp2_index�K�	term2_idx�K u}�(h
�Wire2�h�Kh�Kh�Kh�K u}�(h
�Wire3�h�K h�K h�Kh�Ku}�(h
�Wire4�h�Kh�K h�Kh�K u}�(h
�Wire5�h�Kh�K h�Kh�K u}�(h
�Wire6�h�Kh�Kh�Kh�Ku}�(h
�Wire7�h�Kh�Kh�Kh�Ku}�(h
�Wire8�h�Kh�Kh�Kh�K u}�(h
�Wire9�h�Kh�Kh�Kh�Kue�
comp_index�}�(�resistor�K�voltage_source�K
�current_source�Kuu.
��      }�(�
components�]�(}�(�element��circuit_elements��CircuitElement���)��}�(�name��R1��value�G@�@     �element_type��resistor��nodes�]�(KKeub�	comp_type�h�center�G@h�     G@\      ���rotation�K �shape_points�]�(J����K ��J����J������K K
��K
J������KK ��e�	terminals�]�(J����K ��KK ��e�current_arrows�]�(K$K%e�current��numpy._core.multiarray��scalar����numpy��dtype����f8�����R�(K�<�NNNJ����J����K t�bC      𿔆�R�u}�(hh)��}�(h
�R2�hG@�@     h�resistor�h]�(KK eubhh5hG@s0     G@d�     ��hKZh]�(hhhhheh]�(hheh ]�(K&K'eh"h%h+C      𿔆�R�u}�(hh)��}�(h
�I1�hG?�      h�current_source�h]�(KK eubhhBhG@`      G@e@     ��hKZh]�h]�(hheh ]�(K(K)eh"G?�      u}�(hNh�ground�hG@h�     G@qP     ��hK h]�h]�(J����K ��K
K ��e�	is_ground��h ]�ue�wires�]�(}�(h
�Wire1��comp1_index�K�	term1_idx�K �comp2_index�K �	term2_idx�K u}�(h
�Wire2�hUK hVKhWKhXK u}�(h
�Wire3�hUKhVKhWKhXKu}�(h
�Wire4�hUKhVKhWKhXKue�
comp_index�}�(�resistor�K�voltage_source�K �current_source�Kuu.
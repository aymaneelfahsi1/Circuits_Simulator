��!      }�(�
components�]�(}�(�element��circuit_elements��CircuitElement���)��}�(�name��V1��value�G@      �element_type��voltage_source��nodes�]�(KKeub�	comp_type�h�center�G@u     G@s0     ���rotation�K �shape_points�]��	terminals�]�(K J������K K��e�current_arrows�]�(KNKOe�voltage_arrows�]��current��numpy._core.multiarray��scalar����numpy��dtype����f8�����R�(K�<�NNNJ����J����K t�bC������翔��R�u}�(hh)��}�(h
�V2�hG?�      h�voltage_source�h]�(KKeubhh2hG@z�     G@s     ��hK h]�h]�(hheh]�(KPKQeh]�hh"h(C     �?���R�u}�(hh)��}�(h
�R1�hG@       h�resistor�h]�(KKeubhh@hG@u0     G@f�     ��hKZh]�(J����K ��J����J������K K
��K
J������KK ��eh]�(J����K ��KK ��eh]�(KRKSeh]�hh"h(C������翔��R�u}�(hh)��}�(h
�R2�hG@       h�resistor�h]�(KKeubhhUhG@z�     G@h      ��hKZh]�(hDhEhFhGhHeh]�(hJhKeh]�(KTKUeh]�hh"h(C     �?���R�u}�(hh)��}�(h
�R3�hG@      h�resistor�h]�(KKeubhhchG@��     G@o      ��hKZh]�(hDhEhFhGhHeh]�(hJhKeh]�(KVKWeh]�hh"h(C      �?���R�u}�(hh)��}�(h
�R4�hG@       h�resistor�h]�(K KeubhhqhG@z�     G@z`     ��hK h]�(hDhEhFhGhHeh]�(hJhKeh]�(KXKYeh]�hh"h(C     ࿔��R�u}�(hh)��}�(h
�V3�hG@       h�voltage_source�h]�(KK eubhhhG@x     G@v�     ��hK h]�h]�(hheh]�(KZK[eh]�hh"h(C������߿���R�u}�(hNh�ground�hG@a`     G@x      ��hK h]�h]�(J����K ��K
K ��e�	is_ground��h]�h]�ue�wires�]�(}�(h
�Wire1��comp1_index�K �	term1_idx�K�comp2_index�K�	term2_idx�K u}�(h
�Wire2�h�Kh�Kh�Kh�K u}�(h
�Wire3�h�K h�K h�Kh�Ku}�(h
�Wire4�h�Kh�K h�Kh�Ku}�(h
�Wire5�h�Kh�K h�Kh�K u}�(h
�Wire6�h�Kh�K h�Kh�K u}�(h
�Wire7�h�Kh�Kh�Kh�Ku}�(h
�Wire8�h�Kh�K h�Kh�Ku}�(h
�Wire9�h�Kh�Kh�Kh�Kue�
comp_index�}�(�resistor�K�voltage_source�K�current_source�K uu.
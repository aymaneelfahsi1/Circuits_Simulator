���      }�(�
components�]�(}�(�element��circuit_elements��CircuitElement���)��}�(�name��V1��value�G@@     �element_type��voltage_source��nodes�]�(KK eub�	comp_type�h�center�G@c`     G@rP     ���rotation�KZ�shape_points�]��	terminals�]�(J����K ��KK ��e�current_arrows�]�(MlMme�current��numpy._core.multiarray��scalar����numpy��dtype����f8�����R�(K�<�NNNJ����J����K t�bC      �����R�u}�(hh)��}�(h
�V2�hG@@     h�voltage_source�h]�(KKeubhh0hG@��     G@p�     ��hK h]�h]�(hheh]�(MnMoehh h&C      ࿔��R�u}�(hh)��}�(h
�V3�hG@o@     h�voltage_source�h]�(KKeubhh=hG@�@     G@p�     ��hK h]�h]�(hheh]�(MpMqehh h&C      �?���R�u}�(hh)��}�(h
�R1�hG@�@     h�resistor�h]�(KK eubhhJhG@�H     G@s�     ��hKZh]�(J����K ��J����J������K K
��K
J������KK ��eh]�(hheh]�(MrMsehh h&C      �?���R�u}�(hh)��}�(h
�R2�hG@�@     h�resistor�h]�(KK eubhh\hG@�X     G@t@     ��hKZh]�(hNhOhPhQhReh]�(hheh]�(MtMuehh h&C      �?���R�u}�(hh)��}�(h
�R3�hG@�@     h�resistor�h]�(KKeubhhihG@z�     G@q�     ��hK h]�(hNhOhPhQhReh]�(hheh]�(MvMwehh h&C      ࿔��R�u}�(hh)��}�(h
�R4�hG@�@     h�resistor�h]�(KKeubhhvhG@t�     G@m�     ��hKZh]�(hNhOhPhQhReh]�(hheh]�hh h&C        ���R�u}�(hh)��}�(h
�R5�hG@�@     h�resistor�h]�(KK eubhh�hG@t�     G@s�     ��hKZh]�(hNhOhPhQhReh]�(hheh]�(MxMyehh h&C      �?���R�u}�(hh)��}�(h
�R6�hG@�@     h�resistor�h]�(KK eubhh�hG@o@     G@r      ��hKZh]�(hNhOhPhQhReh]�(hheh]�(MzM{ehh h&C      �?���R�u}�(hNh�ground�hG@d`     G@xp     ��hK h]�h]�(J����K ��K
K ��e�	is_ground��h]�ue�wires�]�(}�(h
�Wire1��comp1_index�K �	term1_idx�K �comp2_index�K�	term2_idx�K u}�(h
�Wire2�h�K h�Kh�Kh�Ku}�(h
�Wire3�h�Kh�K h�Kh�K u}�(h
�Wire4�h�Kh�Kh�Kh�K u}�(h
�Wire5�h�Kh�Kh�Kh�K u}�(h
�Wire6�h�Kh�Kh�Kh�K u}�(h
�Wire7�h�Kh�Kh�Kh�K u}�(h
�Wire8�h�Kh�K h�Kh�K u}�(h
�Wire9�h�Kh�Kh�Kh�K u}�(h
�Wire10�h�Kh�Kh�Kh�Ku}�(h
�Wire11�h�Kh�Kh�Kh�Ku}�(h
�Wire12�h�Kh�Kh�Kh�Ku}�(h
�Wire13�h�K	h�Kh�K h�Kue�
comp_index�}�(�resistor�K�voltage_source�K�current_source�K uu.